* C:\MSimEv_8\Projects\ue4\4_4.sch

* Schematics Version 8.0 - July 1997
* Mon Jul 02 21:50:10 2012



** Analysis setup **
.tran 1us 10ms
.OPTIONS DIGINITSTATE=0
.OP 
.LIB "C:\MSimEv_8\Projects\ue4\4_4.lib"


* From [SCHEMATICS NETLIST] section of msim.ini:
.lib nom.lib

.INC "4_4.net"
.INC "4_4.als"


.probe


.END
