* C:\MSimEv_8\Projects\ue3\1_2.sch

* Schematics Version 8.0 - July 1997
* Sun May 20 19:17:49 2012


.PARAM         Rval=1.1k 

** Analysis setup **
.DC LIN TEMP 0 100 0.1 
+  PARAM Rval LIST 
+ 1089 1100 1111
.OP 
.LIB "C:\MSimEv_8\Projects\ue3\1_2.lib"


* From [SCHEMATICS NETLIST] section of msim.ini:
.lib nom.lib

.INC "1_2.net"
.INC "1_2.als"


.probe


.END
