* Y:\SSIM\UE\REPO\ABGABE4\SIM\2.sch

* Schematics Version 8.0 - July 1997
* Mon Jul 02 22:02:45 2012



** Analysis setup **
.tran 10ns 1.5us
.OPTIONS DIGINITSTATE=2
.OPTIONS DIGIOLVL=1
.OPTIONS DIGMNTYMX=3
.OPTIONS DIGERRDEFAULT=100
.OPTIONS DIGERRLIMIT=100
.STMLIB "2.stl"


* From [SCHEMATICS NETLIST] section of msim.ini:
.lib "nom.lib"
.lib "C:\MSimEv_8\UserLib\SIEMENS.LIB"
.lib "C:\MSimEv_8\UserLib\NAT_SEMI.LIB"
.lib "C:\MSimEv_8\UserLib\mos_int.lib"
.lib "C:\MSimEv_8\UserLib\LIN_TECH.LIB"

.INC "2.net"
.INC "2.als"


.probe


.END
