* Y:\SSIM\UE\Abgabe2\bsp1b.sch

* Schematics Version 8.0 - July 1997
* Thu Mar 22 22:37:15 2012



** Analysis setup **
.OP 


* From [SCHEMATICS NETLIST] section of msim.ini:
.lib nom.lib

.INC "bsp1b.net"
.INC "bsp1b.als"


.probe


.END
