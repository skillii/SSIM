* Y:\SSIM\UE\repo\abgabe3\sim\3_klirr.sch

* Schematics Version 8.0 - July 1997
* Mon May 21 20:36:10 2012



** Analysis setup **
.tran 2ns 0.0035ms 0 0.002us
.OP 


* From [SCHEMATICS NETLIST] section of msim.ini:
.lib "nom.lib"
.lib "C:\MSimEv_8\UserLib\SIEMENS.LIB"
.lib "C:\MSimEv_8\UserLib\NAT_SEMI.LIB"
.lib "C:\MSimEv_8\UserLib\mos_int.lib"
.lib "C:\MSimEv_8\UserLib\LIN_TECH.LIB"

.INC "3_klirr.net"
.INC "3_klirr.als"


.probe


.END
