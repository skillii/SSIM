* Y:\SSIM\UE\REPO\ABGABE4\SIM\1.sch

* Schematics Version 8.0 - July 1997
* Thu Jun 28 12:47:19 2012


.PARAM         BLA=10 

** Analysis setup **
.ac DEC 101 1 100000k
.OP 
.LIB "Y:\SSIM\UE\REPO\ABGABE4\SIM\1.lib"


* From [SCHEMATICS NETLIST] section of msim.ini:
.lib "nom.lib"
.lib "C:\MSimEv_8\UserLib\SIEMENS.LIB"
.lib "C:\MSimEv_8\UserLib\NAT_SEMI.LIB"
.lib "C:\MSimEv_8\UserLib\mos_int.lib"
.lib "C:\MSimEv_8\UserLib\LIN_TECH.LIB"

.INC "1.net"
.INC "1.als"


.probe


.END
