* C:\MSimEv_8\Projects\ue2_ex3\pnp_transfer.sch

* Schematics Version 8.0 - July 1997
* Sat Mar 24 18:06:31 2012



** Analysis setup **
.DC LIN V_V_BE 0 2 0.01 
+  V_V_CE LIST 
+ 10 20 30
.TEMP -10 27 85


* From [SCHEMATICS NETLIST] section of msim.ini:
.lib nom.lib

.INC "3_pnp_transfer.net"
.INC "3_pnp_transfer.als"


.probe


.END
