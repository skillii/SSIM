* C:\MSimEv_8\Projects\ue3\2_2.sch

* Schematics Version 8.0 - July 1997
* Mon May 21 20:08:20 2012


.PARAM         Rval=72 

** Analysis setup **
.ac DEC 1000 10000 1000000
.WCASE AC V([$N_0003]) MAX
+  LIST OUTPUT ALL VARY DEV HI
.TEMP -25 27 100
.LIB "C:\MSimEv_8\Projects\ue3\2_1.lib"
.LIB "C:\MSimEv_8\Projects\ue3\2_2.lib"


* From [SCHEMATICS NETLIST] section of msim.ini:
.lib nom.lib

.INC "2_2.net"
.INC "2_2.als"


.probe


.END
