* C:\MSimEv_8\Projects\ue2_ex3\pmos_output.sch

* Schematics Version 8.0 - July 1997
* Mon Mar 26 20:01:43 2012



** Analysis setup **
.DC LIN V_V_DS 0 20 0.01 
+  V_V_GS LIST 
+ 5 6 7
.TEMP -10 27 85


* From [SCHEMATICS NETLIST] section of msim.ini:
.lib nom.lib

.INC "3_pmos_output.net"
.INC "3_pmos_output.als"


.probe


.END
